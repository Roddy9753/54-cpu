`timescale 1ns / 1ps

//�첽��ȡ���ݣ�ͬ��д��
module DMEM(                    
    input dm_clk,               
    input dm_ena,               
    input dm_r,                 //��ȡʱ����
    input dm_w,                 //д��ʱ����
    input sb_flag,             
    input sh_flag,              
    input sw_flag,             
    input lb_flag,              
    input lh_flag,
    input lbu_flag,     
    input lhu_flag,         
    input lw_flag,           
    input [6:0] dm_addr,        //Ҫ��/д�ĵ�ַ
    input [31:0] dm_data_in,   
    output [31:0] dm_data_out  
    );

reg [31:0] dmem [31:0];//DMEM����

always @(negedge dm_clk) begin
    //ʹ�ܶ˿�����дָ����Ч�Ҷ�ָ����Чʱ������Ĵ�����д������
    if(dm_ena && dm_w &&!dm_r) begin
        if(sb_flag)         //�����SBָ�����Ҫ�Ե�ַ��������
            dmem[dm_addr][7:0] <= dm_data_in[7:0];
        else if(sh_flag)    //�����SHָ���Ҫ�Ե�ַ���Զ�
            dmem[dm_addr >> 1][15:0] <= dm_data_in[15:0];
        else if(sw_flag)    //ʣ�µľ���SWָ���Ҫ�Ե�ַ������
            dmem[dm_addr >> 2] <= dm_data_in;
    end
end

//ʹ�ܶ˿�������ָ����Ч��дָ����Чʱ���Ž���Ӧ��ַ�������ͳ���������Ϊ���迹
assign dm_data_out = (dm_ena && dm_r && !dm_w) ? 
                     (lb_flag ? { {24{dmem[dm_addr][7]}} , dmem[dm_addr][7:0] } : 
                     (lbu_flag ? { 24'h0 , dmem[dm_addr][7:0] } :
                     (lh_flag ? { {16{dmem[dm_addr >> 1][15]}} , dmem[dm_addr >> 1][15:0] } :
                     (lhu_flag ? { 16'h0 , dmem[dm_addr >> 1][15:0] } :
                     (lw_flag ? dmem[dm_addr >> 2]: 32'bz))))) : 32'bz;

endmodule
